//Cache control for FSM & supporting logic. Braydon Burkhardt 2.27.24 rev A

module cache_control (
    input logic clk,
    input logic rst
    
);



endmodule : cache_control
